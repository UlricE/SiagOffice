	
Siag (Scheme In A Grid) %s. No Warranty.	Siag (Scheme In A Grid) %s. Ingen garanti.
File	Arkiv
Edit	Redigera
Block	Block
Format	Format
Data	Data
Plugin	Plugin
Window	F�nster
Plot	Diagram
Tools	Verktyg
Help	Hj�lp
Start another instance of Siag	Starta en ny Siag
Open a Siag document		�ppna ett dokument
Save the contents of the current buffer	Spara det �ppna dokumentet
Preview the contents of the current buffer	F�rhandsgranska det �ppna dokumentet
Print the contents of the current buffer	Skriv ut det �ppna dokumentet
Spelling checker		Stavningskontroll
Cut				Klipp ut
Copy				Kopiera
Paste				Klistra in
Undo				�ngra
Sort ascending			Sortera stigande
Sort descending			Sortera fallande
Plot the contents of the block using lines	Plotta inneh�llet i blocket med hj�lp av linjer
Add the contents of the block	Summera inneh�llet i blocket
Display the Siag online documentation	Visa direkthj�lp f�r Siag
Display the Gnu general public license	Visa Gnu-licensvillkoren
Change the font family	Byt teckensnittsfamilj
Change the font size	Byt teckensnittsstorlek
Change the display style	Byt visningsstil
Change the color	Byt f�rg
Bold text	Fetstil
Italic text	Kursiverat
Left adjusted text		V�nsterjustera
Centered text			Centrera
Right adjusted text		H�gerjustera
Draw grid lines in the block	Rita rutm�nster i blocket
Draw borders around the block	Rita ram runt blocket
Underline the block		Stryk under blocket
Remove grid lines from the block	Ta bort alla linjer fr�n blocket
Select everything		Markera allt
OK				OK
Cancel				Avbryt
File Name:			Filnamn:
Directory:			Katalog:
Select File			V�lj fil
Find				S�k
Extra				Extra
Home				Hem
Examples			Exempel
Family Name			Familjenamn
Size				Storlek
Attributes			Attribut
Borders				Kanter
Adjustment			Justering
Misc				�vrigt
List Selection			Listval
New				Nytt
Open				�ppna
Save				Spara
Save As				Spara som
Preview				F�rhandsgranska
Close				St�ng
Backup Copies			S�kerhetskopior
Settings			Inst�llningar
Margins				Marginaler
Paper Size			Pappersstorlek
Header and Footer		Sidhuvud och sidfot
First Page Number		F�rsta sidnummer
Style				Stil
Foreground Color		F�rgrundsf�rg
Background Color		Bakgrundsf�rg
Enter Date			Mata in datum
Enter Time			Mata in tid
Move Sheet			Flytta ark
Up				Upp
Down				Ned
Edit Applications		Redigera program
Save Applications		Spara program
Applets				Sm�program
Resize				�ndra storlek
Print				Skriv ut
Print Format			Utskriftsformat
Orientation			Orientering
Portrait			St�ende
Landscape			Liggande
Cell Protection			Cellskydd
Respect				Respektera
Ignore				Ignorera
Load External			�ppna externt dokument
Save External			Spara externt dokument
Exit				Avsluta
Undo				�ngra
Delete				Radera
Insert Line			S�tt in rad
Remove Line			Ta bort rad
Insert Column			S�tt in kolumn
Remove Column			Ta bort kolumn
Select All			Markera allt
Select everything		Markera allt
Find				S�k
Find Backward			S�k bak�t
Label				Etikett
SIOD Expression			SIOD-formel
C Expression			C-formel
Guile Expression		Guile-formel
Tcl Expression			Tcl-formel
Change default interpreter	Byt standardtolk
Change Default Interpreter	Byt standardtolk
Other				Annan
Add Property			L�gg till egenskap
Embed Object			B�dda in objekt
Remove Object			Radera objekt
Open Object			�ppna objekt
Save Object			Spara objekt
Set Mark			S�tt m�rke
Set Block			Markera block
Unset Block			Ta bort markering
Copy Block			Kopiera block
Delete Block			Radera block
Fill Block			Fyll block
Smart Fill Block		Fyll block smart
Sort				Sortera
Rows Ascending as Text		Rader stigande som text
Rows Ascending as Numbers	Rader stigande som tal
Rows Descending as Text		Rader fallande som text
Rows Descending as Numbers	Rader fallande som tal
Columns Ascending as Text	Kolumner stigande som text
Columns Ascending as Numbers	Kolumner stigande som tal
Columns Descending as Text	Kolumner fallande som text
Columns Descending as Numbers	Kolumner fallande som tal
Block Sum			Summera blocket
Block Minimum			Minsta v�rde
Block Maximum			St�rsta v�rde
Block Average			Genomsnitt
Borders				Kantlinjer
Grid				Rutm�nster
Underline			Stryk under
None				Inget
Column Width			Kolumnbredd
Set				S�tt
Fit Block			Anpassa till block
Set Default			S�tt standard
Fit Block Width			Anpassa bredd efter block
Row Height			Radh�jd
Fit Block Height		Anpassa h�jd till block
Set Default Format		S�tt standardformat
Cell Format			Cellformat
Block Format			Blockformat
Cell Style			Cellstil
Block Style			Blockstil
Define Style			Definiera stil
Cell Color			Cellf�rg
Block Color			Blockf�rg
Edit Record			Redigera post
Data Entry			Mata in data
Siag-net			Siag-n�tverk
Identify Cell			Identifiera cell
Recalculate			Ber�kna om
Change Buffer			Byt buffer
Delete Buffer			Radera buffer
Split Window			Dela f�nster
Remove Window			Ta bort f�nster
One Window			Ett f�nster
Change Window			Byt f�nster
Add Sheet			L�gg till ark
Remove Sheet			Ta bort ark
Rename Sheet			D�p om ark
Protect Cells			Skydda celler
Remove Protection		Ta bort skydd
Go To				G� till
Beginning of buffer		B�rjan av buffer
End of buffer			Slut av buffer
Top of buffer			Toppen av buffer
Bottom of buffer		Botten av buffer
Grid Lines			Rutm�nster
Show				Visa
Hide				G�m
Reference Style			Referensstil
Disable Helptexts		St�ng av hj�lptexter
Helptexts			Hj�lptexter
Disable				St�ng av
Both				B�da
Save Preferences		Spara inst�llningar
Lines				Linjer
Points				Punkter
Linespoints			Linjer och punkter
Impulses			Streck
Dots				Prickar
Steps				Stegdiagram
Boxes				Staplar
Surface				Ytdiagram
Advanced			Avancerat
Contents			Inneh�ll
Search				S�k
Copying				Upphovsr�tt
About Siag			Om Siag
About Siag...			Om Siag...
About Siag Office...		Om Siag Office...
About Pathetic Writer...	Om Pathetic Writer...
About Egon Animator...		Om Egon Animator...
About Xfiler...			Om Xfiler...
About XedPlus...		Om XedPlus...
About Gvu...			Om Gvu...
Help for Help			Hj�lp f�r hj�lp
Links				L�nkar
Siag Home			Siags hemsida
FTP Directory			FTP-katalog
SIOD Command			SIOD-kommando
C Command			C-kommando
Guile Command			Guile-kommando
Tcl Command			Tcl-kommando
Web Server			Webserver
Mail				Skicka e-post
File Manager			Filhanterare
Form Test			Test av formul�r
Another Form Test		Ett annat test av formul�r
Yet Another Form Test		�nnu ett test av formul�r
Another Form Test Still		Ytterligare ett test av formul�r
Import				Importera
Export				Exportera
Link				L�nka
Move				Flytta
Expression			Formel
Command				Kommando
Sum				Summera
Import Plugin			Importera plugin
Move Plugin			Flytta plugin
Quit				Avsluta
External Program:		Externt program:
Local File			Lokal fil
Compressed File			Komprimerad fil
Archive				Arkiv
Compressed Archive		Komprimerat arkiv
Generic				Allm�nt
Search:				S�k:
Label:				Etikett:
SIOD expression:		SIOD-uttryck:
C expression:			C-uttryck:
Guile expression:		Guile-uttryck:
Tcl expression:			Tcl-uttryck:
New expression interpreter:	Ny formeltolk:
Key				Nyckel
Value				V�rde
Object file:			Objektfil:
Width:				Bredd:
Height:				H�jd:
Bold				Fetstil
Italic				Kursiv
Top				Topp
Bottom				Botten
Left				V�nster
Right				H�ger
Center				Centrera
Expression style:		Uttrycksstil:
Color:				F�rg:
color				f�rg
Black				Svart
Red				R�d
Green				Gr�n
Blue				Bl�
Yellow				Gul
Magenta				Magenta
Cyan				Cyan
White				Vit
Select Plugin:			V�lj plugin:
Change Buffer:			Byt buffer:
Kill Buffer:			Radera buffer:
SIOD command:			SIOD-kommando:
C command:			C-kommando:
Guile command:			Guile-kommando:
Tcl command:			Tcl-kommando:
To:				Till:
Enter user data			Mata in anv�ndardata
First name			F�rnamn
Last name			Efternamn
Address				Adress
Find pattern:			S�k m�nster:
Go to:				G� till:
Pick one:			V�lj en:
Yes				Ja
No				Nej
Replace				Ers�tt
Spell				Stavning
Tab Distance			Tabbavst�nd
Beginning of paragraph		B�rjan av stycke
End of paragraph		Slut av stycke
Line Height			Radh�jd
Segment Format			Segmentformat
Line Format			Radformat
Copy				Kopiera
Use				Anv�nd
Cleanup				St�da
Segment Style			Segmentstil
Line Style			Radstil
Segment Color			Segmentf�rg
Line Color			Radf�rg
About Pathetic Writer		Om Pathetic Writer
Spell Test			Stavningstest
Dump Words			Dumpa ordlista
Default				Standard
Invisible			Osynlig
Integer				Heltal
Scientific			Vetenskaplig
Fixed				Fast
Date				Datum
Time				Tid
Comma				Komma
Percent				Procent
Hex				Hex
Currency			Valuta
User 1				Egen 1
User 2				Egen 2
User 3				Egen 3
User 4				Egen 4
User 5				Egen 5
Header 1			Rubrik 1
Header 2			Rubrik 2
Header 3			Rubrik 3
Header 4			Rubrik 4
Header 5			Rubrik 5
Header 6			Rubrik 6
Title				Titel
Abstract			Utdrag
Preformatted			F�rformaterat
Embed				Inb�dda
Start another instance of Pathetic Writer	Starta en ny Pathetic Writer
Open a Pathetic Writer document		�ppna ett Pathetic Writer-dokument
Display the PW online documentation	Visa direkthj�lpen f�r PW
Underlined text			Understruken text
Superscript			H�jd text
Subscript			S�nkt text
Show Editor			Visa redigerare
Hide Editor			G�m redigerare
Show editor			Visa redigerare
Hide editor			G�m redigerare
Begin Empty Animation		Starta ny animation
Add Object			L�gg till objekt
Line				Linje
Image				Bild
Delete Object			Ta bort objekt
Change Object Type		�ndra objektstyp
Add tick			L�gg till tidpunkt
Delete Tick			Ta bort tidpunkt
Edit Properties			Redigera egenskaper
Set Background			V�lj bakgrund
Timing				Tidsfl�de
Set Geometry			V�lj geometri
Play Animation			Spela upp animation
Box Animation Demo		Demo av boxanimation
Circle Animation Demo		Demo av cirkelanimation
Line Animation Demo		Demo av linjeanimation
Combo Animation Demo		Kombinationsdemo
Box				Rektangel
Circle				Cirkel
Combo				Kombination
About Egon Animator		Om Egon Animator
Start another instance of Egon Animator	Starta en till Egon Animator
Open an Egon Animator document		�ppna ett Egon Animator-dokument
Pop down animation			St�ng animationen
Pause the animation			Pausa animationen
Previous animation frame		Bak�t en bildruta
Play the animation			Spela animationen
Next animation frame			N�sta bildruta
Display the Egon online documentation	Visa direkthj�lpen f�r Egon
Rectangle				Rektangel
Arc					B�ge
Ellipse					Ellips
Pixmap					Pixmap
String					Text
Point					Punkt
Filled Rectangle			Fylld rektangel
Filled Arc				Fylld b�ge
Filled Ellipse				Fylld ellips
Open file				�ppna fil
Save file				Spara fil
Quit animation				Avsluta animationen
Stop animation				Stoppa animationen
Previous frame				Bak�t en bildruta
Next frame				Fram�t en bildruta
Play animation				Spela animationen
Quit Egon				Avsluta Egon
No files found				Inga filer funna
File saved				Fil sparad
This window is too small to split	Detta f�nster �r f�r litet att dela
Couldn't save				Kunde inte spara
Save %s?				Spara %s?
Saved %s				Sparade %s
Saved as %s				Sparad som %s
Loading					Laddar
New file				Ny fil
Load auto startup code?			Ladda automatisk startkod?
Can't open loader file			Kan inte �ppna laddarfil
Parameters:				Parametrar:
External program failed			Externt program misslyckades
Attempt to delete sole ordinary window	Kan inte radera sista f�nstret
No such buffer				Det finns ingen s�dan buffer
Overwrite existing %s?			Skriv �ver befintlig %s?
Can't open saver file			Kan inte �ppna spararfil
Couldn't kill last buffer		Kan inte radera sista buffern
%s command:				%s-kommando:
%s expression:				%s-uttryck:
Already defining kbd macro!		Definierar redan tangentmakro!
Defining kbd macro...			Definierar tangentmakro...
Not defining kbd macro			Definierar inte tangentmakro
Keyboard macro defined			Tangentmakro definierat
Can't execute anonymous macro while defining one	Kan inte utf�ra makro medan det definieras
Input buffer overflow; macro execution terminated	F�r mycket indata; makrodefinition avslutas
Add Tick				L�gg till tidpunkt
Add Line				L�gg till linje
Add Rectangle				L�gg till rektangel
Add Arc					L�gg till b�ge
Add Ellipse				L�gg till ellips
Add Image				L�gg till bildfil
Add String				L�gg till text
Add Point				L�gg till punkt
Add Filled Rectangle			L�gg till fylld rektangel
Add Filled Ellipse			L�gg till fylld ellips
Add Filled Arc				L�gg till fylld b�ge
Sheet %d				Ark %d
Section %d				Avsnitt %d
Alert					Varning
All files (*)				Alla filer (*)
Change %s:				�ndra %s:
Duration				Varaktighet
ERROR					FEL
Font					Typsnitt
LABEL					ETIKETT
EMPTY					TOM
No object selected			Inget objekt valt
No warranty				Ingen garanti
Object type:				Objekttyp:
Previewer				F�rhandsgranskare
Print Command				Utskriftskommando
Save %s ?				Spara %s ?
Saving					Sparar
Style %s changed			Stil %s �ndrad
This command does nothing		Detta kommando g�r ingenting
Time Difference				Tidsskillnad
Time:					Tid:
black					svart
blue					bl�
cyan					cyan
done.					klart.
green					gr�n
magenta					magenta
white					vit
yellow					gul
yes					ja
Directories				Kataloger
Files					Filer
Top:					Topp:
Bottom:					Botten:
Left:					V�nster:
Right:					H�ger:
Header:					Sidhuvud:
Footer:					Sidfot:
Size:					Storlek:
Respect protection			Respektera cellskydd
Date:					Datum:
Type:					Typ:
Orientation:				Orientering:
Logarithmic X axis			Logaritmisk X-axel
Logarithmic Y axis			Logaritmisk Y-axel
Has ticks				Har ticks
Has titles				Har titlar
Parametric				Parametrisk
Integration				Integrering
Printer					Skrivare
Editor					Editor
Help browser				Hj�lpl�sare
File manager				Filhanterare
Header on first page			Sidhuvud p� f�rsta sidan
Name:					Namn:
Special Char				Specialtecken
Code:					Kod:
Word:					Ord:
Tab distance:				Tabbavst�nd:
First page number:			F�rsta sidnummer:
Height:					H�jd:
Can't make postscript			Kan inte skapa postscript
Objects					Objekt
Ticks					Tidpunkter
Properties				Egenskaper
None selected				Inget valt
Width					Bredd
Height					H�jd
Visible					Synlig
[%s at %d] [size = %dx%d] [duration=%d delta=%d]	[%s vid %d] [storlek = %dx%d] [varaktighet=%d avst�nd=%d]
Line in buffer				Rad i buffern
Line:					Rad:
Insert					Infoga
Save Selection				Spara markerat
Print Selection				Skriv ut markerat
Shift Selection Right			Skifta markerat �t h�ger
Shift Selection Left			Skifta markerat �t v�nster
Jump					Hoppa
Begin					Start
End					Slut
Selection Start				Start av markering
Selection End				Slut av markering
Search Selection			S�k markerat
Replace Selection			Ers�tt markerat
Find Bracket				Finn parentes
Check Brackets				Kontrollera parenteser
Options					Inst�llningar
Call Sed				Anropa Sed
About					Om
Commands				Kommandon
New Xedplus				Ny Xedplus
Pipes					R�rledningar
Pipe					R�rledning
-Insert-				-Infoga-
-Overwrite-				-Skriv �ver-
Start another editor			Starta ny editor
Open a text file			�ppna textfil
Save the file				Spara filen
Print the file				Skriv ut filen
Display the online documentation	Visa direkthj�lp
no file yet				�nnu ingen fil
Line number?				Radnummer?
Start at:				B�rja vid:
Cursor position				Ins�ttningspunkt
Textbeginning				Textstart
Textending				Textslut
Direction:				Riktning:
Forward					Fram�t
Backward				Bak�t
Search for:				Leta efter:
Replace with:				Ers�tt med:
Replace veto				Ers�tt fr�ga
Replace all				Ers�tt alla
Wrap mode:				Radbrytningss�tt:
Never					Aldrig
Word					Ord
Tab size:				Tabbavst�nd
Autoindent:				Autoindentera:
Autofill:				Autofyll:
Perform a stream editor command (sed)	Utf�r ett str�meditorkommando (sed)
Command:				Kommando:
Do it					Utf�r
Do it Selection				Utf�r p� markering
Undo it					�ngra
Perform a User command			Utf�r ett anv�ndarkommando
Perform a User pipe			Utf�r ett r�rledningskommando
New...					Nytt...
Move...					Flytta...
Copy...					Kopiera...
Link...					L�nka...
Select...				Markera...
Select all				Markera allt
Deselect all				Avmarkera allt
Folder					Katalog
Go to...				G� till...
Empty					T�m
View					Visa
Tree					Tr�d
Icons					Ikoner
Text					Text
Sort by name				Sortera efter namn
Sort by size				Sortera efter storlek
Sort by date				Sortera efter datum
Hide folders				G�m kataloger
Mix folders/files			Blanda kataloger/filer
Show hidden files			Visa g�mda filer
Close window				St�ng f�nstret
Go to home directory			G� till hemkatalogen
Go up one directory			G� upp en katalog
Create folder				Skapa katalog
Open command window			�ppna kommandof�nster
Change view mode			�ndra visningss�tt
Change sort mode			�ndra sorteringss�tt
Text editor				Texteditor
Find file				S�k efter fil
Create file:				Skapa fil:
Filename pattern:			Filnamnsm�nster:
Add					L�gg till
Remove					Ta bort
Create folder:				Skapa katalog:
Go to folder:				G� till katalog:
Clear					Rensa
Copy to:				Kopiera till:
Move to:				Flytta till:
Link to:				L�nka till:
Command Window				Kommandof�nster
Information...				Information...
Name					Namn
Length					L�ngd
Owner					�gare
Group					Grupp
Access Permissions			R�ttigheter
Type					Typ
Symbolic Link To			Symbolisk l�nk till
Last Modification			Sista inneh�lls�ndring
Last Status Change			Sista status�ndring
Permissions...				R�ttigheter...
Changing access permissions for %s	�ndrar r�ttigheter f�r %s
Others					�vriga
Restore					�terst�ll
Open With...				�ppna med...
Open with:				�ppna med:
Redo					Igen
Stop					Stopp
Open...					�ppna...
Reopen					�ppna igen
Print...				Skriv ut...
Print marked pages...			Skriv ut markerade sidor...
Save marked pages...			Spara markerade sidor...
Page					Sida
Next					N�sta
Redisplay				Visa igen
Previous				F�reg�ende
Mark					Markera
Unmark					Ta bort markering
Magstep					Storlek
Upside-down				Upp och ner
Seascape				Liggande upp och ner
Swap Landscape				Omv�nt liggande
Help...					Hj�lp...
Copyright...				Copyright...
Open a PostScript file			�ppna en Postscriptfil
Save the marked pages			Spara de markerade sidorna
Print the marked pages			Skriv ut de markerade sidorna
Previous page				Bak�t en sida
Next page				Fram�t en sida
Center page				Centrera sidan
Increase magstep			St�rre
Decrease magstep			Mindre
Display online help			Visa direkthj�lp
Display copyright information		Visa copyrightinformation
Printer Name:				Skrivarens namn:
Okay					OK
Unsaved Changes!			�ndringar �r inte sparade!
File has been modified by someone else!	Filen har �ndrats av n�gon annan!
Cannot create backup file!		Kan inte skapa s�kerhetskopia!
Cannot open file for reading!		Kan inte �ppna filen f�r l�sning!
File does not exist and directory is write protected!	Filen finns inte och katalogen �r skrivskyddad!
File opened READ ONLY			Filen �ppnad SKRIVSKYDDAD
Cannot open file!			Kan inte �ppna filen!
Cannot save file!			Kan inte spara filen!
Cannot create file!			Kan inte skapa filen!
Error in Print Command String		Fel i skrivarkommando
Don't know how to handle this drop!	Kan inte hantera detta sl�pp!
Update icons				Uppdatera ikoner
Which format?				Vilket format?
Warning!				Varning!
Warning					Varning
Toggle overwrite/insert			V�xla mellan �verskrivning och ins�ttning
This program is part of Siag Office,\nan effort to create a full-featured, free\noffice package for Unix and X.		Detta program �r en del av Siag Office,\nett projekt f�r att skapa ett komplett\nofficepaket f�r Unix och X.
The interactive text editor for X	Den interaktiva texteditorn f�r X
Authors:				Programmerare:
Part of Siag Office			Del av Siag Office
A spreadsheet for X			Ett kalkylprogram f�r X
A word processor for X			Ett ordbehandlingsprogram f�r X
An animation program for X		Ett animeringsprogram f�r X
A file manager for X			En filhanterare f�r X
A postscript viewer for X		En postscriptvisare f�r X
Environment				Milj�
Custom					Special
Defaults				Standard
Calculator				Kalkylator
Leftline the block			Linjer till v�nster
Rightline the block			Linjer till h�ger
Clear Background			T�m bakgrund
Set Gradient				S�tt gradient
Clear Gradient				Ta bort gradient
Strikethrough				Genomstruken
Full adjusted text			Fulljusterad text
Close Buffer				St�ng buffer
File saved via external program		Filen sparades av externt program
Save %s before checking spelling?	Spara %s f�re stavningskontroll?
Edit Tabs				Redigera tabbar
Theme					Tema
Restart to activate theme		Starta om f�r att aktivera tema
No theme selected			Inget tema valt
Select					V�lj
